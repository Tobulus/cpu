`ifndef mem_acc_vh
`define mem_acc_vh
    localparam MEM_NOP   = 2'b00;
    localparam MEM_READ  = 2'b01;
    localparam MEM_WRITE = 2'b10;
`endif
