`ifndef cmp_res_vh
`define cmp_res_vh
    localparam CMP_EQ = 0;
    localparam CMP_RA_GT = -1;
    localparam CMP_RB_GT = 1;
`endif
